��/  K��@AZ�����"SƤ`��g�o[j#ƽ�n-1��͈�P�Ǜ�*e�c�1��E#nT-�}�Ւ���݆C��=��a��	z>���:Аͭ���0/6q���qrP�@�u���m��U�*�VJ��$+ߴ���V��$b�]_�;R�߭"""�k�{��1����]U�h6O��ȫ���� �����>��zܭQe�^V����R�0��:�@�x�CL[�������ě�o�E�!��*���K��S�nhצr-�Q.��vL��s��T@�t�c1��!V�7�t�Y0��Z��cW0�R��Mm����)
�r�&��MR�Ѧ�	�����.������CC��Q��n$Ӏl!�#*&�E6��1�6Jx�B�m��[�j?��^���<?��>f#-|�-��oB���ޕ�{��ѩ�ƪD��s�xsٸ�Z�0��I�"ㅊ�L�O�D���d�\�Tc���8�^pr�m��4[����,���Kk���=g�
9g���������X��⼑gC� �h������0�i��<t7�LO�6h��;��7,݄�"^4>�1���v�X.�v�$�9�9a�kd��16@%�}�zer�`n��Ą�O�̭u��|�!��Nk���Gϒ!�}��U�7�]�{�mØ�vС�7A�
�s�nk7r&yp"�Os����%%,�O��}+.��I�[�OQ9�soP���:*l���F���Uti�|t��̱Lzࡂ��,�"�w)/�O6T�o�����W\�RI�gZGZ��W��L�W��.,� �Q�����|���]܁4��$ �k��WZzy��N�X�F�0�3��HL��*�U6K4��̕��	ۣ����CKwtR���X��[�4;���#�Nm�E�;�e�R��(+�B���X�1�͂��>���iI�<���r��u��͘{&f����-?6t�<V|r%S-��0���Y���[� i���}l��⚮R�dz�������	�Q�l_Fʵ��@Z�r�Pj���I�ؚ^ᇌߧP.�Z=��#�y���g�!1
���Ɇ��F1 J�S��V�e�W����7 ���hoM�F/�r�w6��w�4g��p��]��||�^x�-JPEp:�+��*�a�ٲb�uR�/lq6D���]+�5�bok��.{2��JS���U � L�%s!��5���M�ڌb��w7�MX�e5���#���(W�2Z���S����<���qs;�{���g��k��M�?��g����pj��æ�5�Qv�*�5+�+���)�1�6�[�ݽ˓�%.���瀂eS�����n��6�a�>
=I|�j}�� ���3ǣ�> �z�����+g���=?��S�cB���(��%L	���`dƞ�4]=��Q��:�*p}�w,MSTZ��AC�i��ʛ���Z�­.&#[�_e�������Zֺ��I|�?�'FfB�W�ԧF�����hʘkl��J/�I�	L�!�ud孝(	]�u��s2���s��4/���g��n"=��.�z�p1�2�e���t��ω8��Ji���1��H5���']�
:ب�a1�.-��[o��8i]���z`�(J���a�^;_�];j�L�����.�
�V!�m*��]c�����z:^h��+�qy�Zqs�Y���>�J��~�����`aWR�����m�����Y�(��
�fF���D��ӓdjUգ����T��ey,Z�n6�E�$3-�$�Yz�[�f��
hL娡Y�+{��,3�<M�t�����=�#H}�k:Q��{�F���tk�E�&{�c�-�G�I�vV抜O�ru2��޷<�O@���%?��T���.��u����ۋr�j����[���\;2��kh��| ���vǃ(PLp��;ߝ����DB4�������i�#����t��f�;��?R�gv����V�#�c�s������e>j���9h�+��q)�=>	
L��'�%щQ.Eq����g�<kSӃfKr�h{�c��9��hqK����GW*R��l���~�WzWPs]�g8Z�fZ$�k�G��y�/u���å� P��3��Dy���3�<�>�z�b�J٘~��3���ީh\y��f��%PO�+[�������D�-�G�%7rz�Z��rw�	,
�*
�*L��0�`�BunQ|�_�y�ޣ�$�̖nH��(�A)�"ھ�ʲ�I�v�C�|G�niY@��<�0^=����C(�z�t�v aԩ�0N3dw���2}m�4�?�N�td�f�)���Mq��*%��w��z������� m
K?v)��׎w��׼S����0C�+����L��1/�R2�f�6� |�ȪA��\�u��:Y������&J�]���?7�CP�*�',u��/�I��$U��1�*K�oTr��6��-���Fś�g���!���"{����QH���na��C��Fa\���n��f`PˁȀ^
gwR۲�f88q"�a�����0zm����[<�c�bA���G ia�.�64���(��k���]o��=�+ ��m���$��u#Iֽ�
����l$�Kk���]��ٵ�Iψ��-��1`u�o�T�h��䳸���뺛oq�([�C��_+�+٠a�w|Vϕ�NI��H��	Fpw�
;��֊h�~�4gǘp��P�`0�r`^�" t`-cٷDځH��}`ji(��n�)/�����Q_����g�{t��9�
`�Y+߻^���9!�%z��� �i��~�\_�6h����i1z|���V�.�:�"�G����\>q�ˎ��<5N��p(��� ��Ϲ�����L���u�=#g$��wq�[�ۣ��	�� #����5yu5��Z���5����v�&������{q�n�i���y��$�D,��))�}�-��_w�h����o��]���t�jQ&�_�� ��EvKO86G3:f���	�{uL4�36&{�w�2�&��9�Y0�)��$/�����;�=f�O�v��C�Ӛ$��8��>��G>��Ebf��Oz��P?�].�]���_�?������|4��)X�lVҰ�a��%�9#i׶�ﵮ�7�� ��`��+C��<�[/#���,���8�|�7k��H����5ʺ$��2v�HE�4�[����J�1���ّ:��rp� ���U<��L�B�Հ���h�C�OZ�!���J���!=Q���.MiMo��$�����o�?By��E��*Ћ����ñ�4Tc +ȳ�	k*�5�Ӏ��˕D��f��&p�\�>Xm.�=�._
����ts�6��I^�мO�Fsj�/rM
)b�׽%`�\��pʱm�[�Yz���/|1���q�߼?�%�ٴğ��>�]E*FF��N�Ϋ:m���/u6��CL��z��i6��"���;0���KtYq(/��op������u�ɵq���HE�˂���P�g'|ϳ;�i�������Z�o��d���&�w�������77��{�+]x�eQ�͟�	�4<WW��_��J�K�����8��*�
����m�5C3�{�A���:�0YB���\2��|+7�"�Tz|��'�c���nuU�K]���I裱�'��o��mlU0�ϱ���!CJ>����i���d��-H�=�>�;/%;��C��DO��k_�!0ީ��_Ε".�k�?]����T�,�Yi#j|���η��-�xa�XtЅϬ�٥ӧ�����m�ͩ����# �>�_ۦ��1�)�$���h�U�I$�;W��"��b��K� Tz>�bnO�zmT`0Sb7P�镳��Z��႒��	�hjݓ�`r�P9�7A��G^n|�9o���E���j[�$�p��K+#Xĥ/�f2�+$Pz��2(4恱)��|0�O�hѯ1�p�Hiv���J�Q.o��wB���N��H�`Q�E�� r�]w��b;�:�g�;b��キ�aR޽Ng|�0�v��\�
$Y8M�C3��6����;���[xŜN�pTr��W�skR^V������"��"C�h��;C�e"O�78m��l�3ԓ�@l���hln�O����V���"G��'t�v�\�Z2�i8�9�0�(\��2Yp_�[gg�G+��X���msW�7�u�?�jl��	�Kv��q�������F5� h��#��~u��4`���-�]!���Sa$x�c�����I�
�4u�S�q3���_ #;��{�Ӱ;�)�(s�1`�t��^��'�MO���I�d倃=H{ޭ��G�0��Ds5�܈V��{{�}~l�Gy�oNp�k.�!�m�l|j5��OS{cQ͟#(w(�h˵0��Ϲ
S�[Ԕ�'����!��a��w�s)W�t����d.��ZS:�Tx,@\���o��דM��Ȋ-���^�dZd��Y=%2�^S���Ô��~-ס!�eG���H�:���g��j�]����bI��@�R���AXY?��~�ҹ`T�r���վ��0��*����Qw~Wk�QT�a���3%�D�bifR�-F��Y%�oX��O֨�\T&i|X�_k�v�q�*���?Kv�����Y�**���Vz[[��A���4P\�vkD��q��ŹҺjÄ9f݋��&4�bʉO+Q�����ߛ�����Ck�2X��kR�ع�/Z9J_j�����a{a41{+J�[��@-x�_ 6��d.m�~����1Jz�~RYv�O!���쩀 �>r5J�,�ĝ�7�zx(-B��=֟��jvh�D�,A�7�)��B2�z�����xu�8I�o�}�\������L�W0�Z����iF7�!�]�2�F����������/�����hGa��џ;���m��)WM�����@�=���6zt��+q۵<�����E�W;�س���E�ayq��vAq\�v��=��>~/L�!�!+˅B��^�X�?d�&H�6�t��xe9�"��;Ɨ����je���� T���,mM��jc	L�U�b��X��c����a��$qOwuA�ΎPgu�c<vY>��r����q��3ds�5�Fd�����q)ҴsT��L�J\�d�bc��ؒ��(�H=Z�cu�jP�0:MMIXp������09��9Xra� d�}�O$E�	�H�V�Aج2�F�|/6�+S��K{*��1)PT	(B��`��H��x�'�|���O���s���o��A�Q����.O����(��|Ys���Y
��H5��^R�Xg�7e���m�B�%�L�(F�;QA��t��5A.���|6A���^:?�IU��n�L��)����CN�v�iL*,߈�QI����zƅ�K-��c�J��oe�M^��{�K5D�e�~���9���f0�v4��nc������}�L���Ks��D-�Pzj@�ŧى��